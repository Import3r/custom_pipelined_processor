module testSub();
reg [7:0] x,y;
wire [3:0] st;
wire [7:0] res;
initial begin
x<=8'b00000001; y<=8'b00000001; //0
#25 x<=8'b00000100; y<=8'b00000001; //3
#25 x<=8'b01111111; y<=8'b00000001; //126
#25 x<=8'b01111111; y<=8'b00000111;//120
#25 x<=8'b01101011; y<=8'b01000000;//43
#25 x<=8'b10000000; y<=8'b00000000;//-128
#25 x<=8'b01111000; y<=8'b11110111; //120-(-9) -> overflow
#25 x<=8'b01111000; y<=8'b00001001;//120-9 
#25 $finish;
end
sub s1(x,y,res,st);
endmodule