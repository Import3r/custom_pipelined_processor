module instructionMemory(instruction, PC);

	integer j;
	input [31:0]PC;
	output [31:0]instruction;
	reg [7:0] mem [16383:0];
	wire [31:0]instruction;
	initial begin
			// SOME softwares would have a 5000 limit on for loop.
			// You can break this into multiple loops or initialize several locations in parallel
			/*for (j = 0; j<4999; j = j + 1)//16k
				begin
					mem[j] <= 8'b0;
				end		
			for (j = 5000; j<10000; j = j + 1)//16k
				begin
					mem[j] <= 8'b0;
				end				
			for (j = 10001; j<15000; j = j + 1)//16k
				begin
					mem[j] <= 8'b0;
				end
			for (j = 15001; j<16384; j = j + 1)//16k
				begin
					mem[j] <= 8'b0;
				end*/
				
			// ******************************************************	
			///Test Case 1: Load Operations 
			// ****************************************************** 
			//lw $t0,0($0)
			//lw $t1,4($0)
			//lw $t2,8($0)
			//lw $t3,12($0)
			//lw $t4,16($0)
			//lw $t5,20($0)
			//lw $t6,24($0)
			//lw $t7,28($0)
			
				
			mem[100] <= 'h48;
			mem[101] <= 'h08;
			mem[102] <= 'h00;
			mem[103] <= 'h00;
			
			mem[104] <= 'h48;
			mem[105] <= 'h09;
			mem[106] <= 'h00;
			mem[107] <= 'h04;
			
			mem[108] <= 'h48;
			mem[109] <= 'h0a;
			mem[110] <= 'h00;
			mem[111] <= 'h08;
			
			mem[112] <= 'h48;
			mem[113] <= 'h0b;
			mem[114] <= 'h00;
			mem[115] <= 'h0c;
			
			mem[116] <= 'h48;
			mem[117] <= 'h0c;
			mem[118] <= 'h00;
			mem[119] <= 'h10;
			
			mem[120] <= 'h48;
			mem[121] <= 'h0d;
			mem[122] <= 'h00;
			mem[123] <= 'h14;
			
			mem[124] <= 'h48;
			mem[125] <= 'h0e;
			mem[126] <= 'h00;
			mem[127] <= 'h18;
			
			mem[128] <= 'h48;
			mem[129] <= 'h0f;
			mem[130] <= 'h00;
			mem[131] <= 'h1c;
			
			// ******************************************************	
			///Test Case 2: Arithematic operations - No Forwarding
			// ****************************************************** 
			//addi $s1,$0,5
			//addi $s2,$0,10
			//addi $s3,$0,3
			//addi $s4,$0,2			
			//add  $s5,$s1,$s2
			//sub  $s6,$s1,$s3
			mem[200] <= 'h24;
			mem[201] <= 'h13;
			mem[202] <= 'h00;
			mem[203] <= 'h05;
			
			mem[204] <= 'h24;
			mem[205] <= 'h14;
			mem[206] <= 'h00;
			mem[207] <= 'h0a;
			
			mem[208] <= 'h24;
			mem[209] <= 'h15;
			mem[210] <= 'h00;
			mem[211] <= 'h03;
			
			mem[212] <= 'h24;
			mem[213] <= 'h16;
			mem[214] <= 'h00;
			mem[215] <= 'h02;
			
			mem[216] <= 'h0e;
			mem[217] <= 'h74;
			mem[218] <= 'hb8;
			mem[219] <= 'h20;
			/*Habed Statrt
			mem[212] <= 'hAC;
			mem[213] <= 'h13;
			mem[214] <= 'h00;
			mem[215] <= 'h00;
			
			mem[216] <= 'h48;
			mem[217] <= 'h16;
			mem[218] <= 'h00;
			mem[219] <= 'h00;
			//Habed End*/
			mem[220] <= 'h0e;
			mem[221] <= 'h75;
			mem[222] <= 'hc0;
			mem[223] <= 'h24;
			//Habed
			//addi
			mem[224] <= 'h14;
			mem[225] <= 'h00;
			mem[226] <= 'hFF;
			mem[227] <= 'hE0;
			//beq
			mem[228] <= 8'b00010101;
			mem[229] <= 8'b00101010;
			mem[230] <= 8'b11111111;
			mem[231] <= 8'b11111000;
			//SRL
			mem[232] <= 'h0c;
			mem[233] <= 'h09;
			mem[234] <= 'h88;
			mem[235] <= 'h42;
					//lui
			mem[236] <= 'h3c;
			mem[237] <= 'h0f;
			mem[238] <= 'h00;
			mem[239] <= 'h0a;
			//sw
			mem[240] <= 'had;
			mem[241] <= 'h2a;
			mem[242] <= 'h00;
			mem[243] <= 'h02;
			//lw
			mem[244] <= 'h48;
			mem[245] <= 'h16;
			mem[246] <= 'h00;
			mem[247] <= 'h07;
			//Jr t8 = 232
			//0c090008
			/*mem[296] <= 'h0c;
			mem[297] <= 'h09;
			mem[298] <= 'h00;
			mem[299] <= 'h08;*/
			//JAL 1c00003a
			/*mem[296] <= 'h1c;
			mem[297] <= 'h00;
			mem[298] <= 'h00;
			mem[299] <= 'h3a;*/
			//j 232
			/*mem[296] <= 'h08;
			mem[297] <= 'h00;
			mem[298] <= 'h00;
			mem[299] <= 'h3A;			*/
		//swn 4 0x0C0A4813
			mem[292] <= 'h0C;
			mem[293] <= 'h0A;
			mem[294] <= 'h48;
			mem[295] <= 'h13;	
	//lwn 4 0x0C0F4821
			mem[296] <= 'h0C;
			mem[297] <= 'h0F;
			mem[298] <= 'h48;
			mem[299] <= 'h21;
			// ******************************************************	
			///Test Case 3: Logical Operations - No Forwarding
			// ****************************************************** 
			//addi $s1,$0,15
			//addi $s2,$0,10
			//addi $s3,$0,3
			//addi $s4,$0,2			
			//and  $s5,$s1,$s2
			//or   $s6,$s2,$s3
			mem[300] <= 'h24;
			mem[301] <= 'h13;
			mem[302] <= 'h00;
			mem[303] <= 'h0F;
			
			mem[304] <= 'h24;
			mem[305] <= 'h14;
			mem[306] <= 'h00;
			mem[307] <= 'h0a;
			
			mem[308] <= 'h24;
			mem[309] <= 'h15;
			mem[310] <= 'h00;
			mem[311] <= 'h03;
			
			mem[312] <= 'h24;
			mem[313] <= 'h16;
			mem[314] <= 'h00;
			mem[315] <= 'h02;
			
			mem[316] <= 'h0e;
			mem[317] <= 'h74;
			mem[318] <= 'hb8;
			mem[319] <= 'h14;
			
			mem[320] <= 'h0e;
			mem[321] <= 'h95;
			mem[322] <= 'hc0;
			mem[323] <= 'h25;

			// ******************************************************	
			///Test Case 4: Store Operation
			// ****************************************************** 
			//addi $s1,$0,15
			//addi $s2,$0,10
			//addi $s3,$0,3
			//sw   $s1,100($0)			
			//addi $s1,$0,0
			//addi $s2,$0,10			
			//lw   $s3,100($0)						

			mem[400] <= 'h24;
			mem[401] <= 'h13;
			mem[402] <= 'h00;
			mem[403] <= 'h0f;
			
			mem[404] <= 'h24;
			mem[405] <= 'h14;
			mem[406] <= 'h00;
			mem[407] <= 'h0a;
			
			mem[408] <= 'h24;
			mem[409] <= 'h15;
			mem[410] <= 'h00;
			mem[411] <= 'h03;
			
			mem[412] <= 'hac;
			mem[413] <= 'h13;
			mem[414] <= 'h00;
			mem[415] <= 'h64;
			
			mem[416] <= 'h24;
			mem[417] <= 'h13;
			mem[418] <= 'h00;
			mem[419] <= 'h00;
			
			mem[420] <= 'h24;
			mem[421] <= 'h14;
			mem[422] <= 'h00;
			mem[423] <= 'h0a;
			
			mem[424] <= 'h48;
			mem[425] <= 'h15;
			mem[426] <= 'h00;
			mem[427] <= 'h64;			
			
			// ******************************************************	
			///Test Case 5: Branch Equal - Not Taken
			// ****************************************************** 
			//addi $s1,$0,15
			//addi $s2,$0,10
			//addi $s3,$0,3
			//addi $s4,$0,2			
			//beq  $s1,$s2,-5
			//addi $s1,$0,30
			//addi $s2,$0,20
			//addi $s3,$0,6
			//addi $s3,$0,6
			//addi $s3,$0,6						
		
			mem[500] <= 'h24;
			mem[501] <= 'h13;
			mem[502] <= 'h00;
			mem[503] <= 'h0f;
			
			mem[504] <= 'h24;
			mem[505] <= 'h14;
			mem[506] <= 'h00;
			mem[507] <= 'h0a;
					
			mem[508] <= 'h24;
			mem[509] <= 'h15;
			mem[510] <= 'h00;
			mem[511] <= 'h03;
					
			mem[512] <= 'h24;
			mem[513] <= 'h16;
			mem[514] <= 'h00;
			mem[515] <= 'h02;
			
			// BEQ
			mem[516] <= 'h16;
			mem[517] <= 'h74;
			mem[518] <= 'hff;
			mem[519] <= 'hfb;
			
			mem[520] <= 'h24;
			mem[521] <= 'h13;
			mem[522] <= 'h00;
			mem[523] <= 'h1e;
					
			mem[524] <= 'h24;
			mem[525] <= 'h14;
			mem[526] <= 'h00;
			mem[527] <= 'h14;
					
			mem[528] <= 'h24;
			mem[529] <= 'h15;
			mem[530] <= 'h00;
			mem[531] <= 'h06;			
			
			mem[532] <= 'h24;
			mem[533] <= 'h15;
			mem[534] <= 'h00;
			mem[535] <= 'h06;
					
			mem[536] <= 'h24;
			mem[537] <= 'h15;
			mem[538] <= 'h00;
			mem[539] <= 'h06;	
		

			// ******************************************************	
			///Test Case 6: ALU-ALU FWD 
			// ****************************************************** 
			//addi $s1,$0,15
			//addi $s2,$0,10
			//addi $s3,$0,3
			//add  $s4,$s1,$s2			
			//add  $s5,$s4,$s3
			
			mem[600] <= 'h24;
			mem[601] <= 'h13;
			mem[602] <= 'h00;
			mem[603] <= 'h0f;
			
			mem[604] <= 'h24;
			mem[605] <= 'h14;
			mem[606] <= 'h00;
			mem[607] <= 'h0a;
			
			mem[608] <= 'h24;
			mem[609] <= 'h15;
			mem[610] <= 'h00;
			mem[611] <= 'h03;
			
			mem[612] <= 'h0e;
			mem[613] <= 'h74;
			mem[614] <= 'hb0;
			mem[615] <= 'h20;
			
			mem[616] <= 'h0e;
			mem[617] <= 'hd5;
			mem[618] <= 'hb8;
			mem[619] <= 'h20;
//OUR-TEST-CASE
// lw $t0 0($0)
mem[700] <= 8'b01001000;
mem[701] <= 8'b00001000;
mem[702] <= 8'b00000000;
mem[703] <= 8'b00000000;

// addi $t0 $t0 2
mem[704] <= 8'b00100101;
mem[705] <= 8'b00001000;
mem[706] <= 8'b00000000;
mem[707] <= 8'b00000010;

// andi $t0 $t0 2
mem[708] <= 8'b00110001;
mem[709] <= 8'b00001000;
mem[710] <= 8'b00000000;
mem[711] <= 8'b00000010;

// sll $t0 $t0 2
mem[712] <= 8'b00001100;
mem[713] <= 8'b00001000;
mem[714] <= 8'b01000000;
mem[715] <= 8'b10000000;

// srl $t0 $t0 1
mem[716] <= 8'b00001100;
mem[717] <= 8'b00001000;
mem[718] <= 8'b01000000;
mem[719] <= 8'b01000010;

// nor $t0 $t0 $s0
mem[720] <= 8'b00001101;
mem[721] <= 8'b00010010;
mem[722] <= 8'b01000000;
mem[723] <= 8'b00100111;

// sw $t0 0($0)
mem[724] <= 8'b10101100;
mem[725] <= 8'b00001000;
mem[726] <= 8'b00000000;
mem[727] <= 8'b00000000;

// addi $t1 $0 6
mem[728] <= 8'b00100100;
mem[729] <= 8'b00001001;
mem[730] <= 8'b00000000;
mem[731] <= 8'b00000110;

// addi $t2 $0 6
mem[732] <= 8'b00100100;
mem[733] <= 8'b00001010;
mem[734] <= 8'b00000000;
mem[735] <= 8'b00000110;

// sub $t1 $t1 $t2
mem[736] <= 8'b00001101;
mem[737] <= 8'b00101010;
mem[738] <= 8'b01001000;
mem[739] <= 8'b00100100;

// lwn $t2 $0 $t1
mem[740] <= 8'b00001100;
mem[741] <= 8'b00001010;
mem[742] <= 8'b01001000;
mem[743] <= 8'b00100001;


// addi $t3 $t2 16
mem[744] <= 8'b00100101;
mem[745] <= 8'b01001011;
mem[746] <= 8'b00000000;
mem[747] <= 8'b00010000;

// addi $t1 $0 2
mem[748] <= 8'b00100100;
mem[749] <= 8'b00001001;
mem[750] <= 8'b00000000;
mem[751] <= 8'b00000010;

// addi $t2 $0 2
mem[752] <= 8'b00100100;
mem[753] <= 8'b00001010;
mem[754] <= 8'b00000000;
mem[755] <= 8'b00000010;

// swn $t3 $t1 $t2
mem[756] <= 8'b00001101;
mem[757] <= 8'b01001011;
mem[758] <= 8'b01001000;
mem[759] <= 8'b00010011;

// lbu $t4 7($0)
mem[760] <= 8'b10001000;
mem[761] <= 8'b00001100;
mem[762] <= 8'b00000000;
mem[763] <= 8'b00000111;

// add $t0 $t1 $t2
mem[764] <= 8'b00001101;
mem[765] <= 8'b00101010;
mem[766] <= 8'b01000000;
mem[767] <= 8'b00100000;

// or $t0 $t0 $t1
mem[768] <= 8'b00001101;
mem[769] <= 8'b00001001;
mem[770] <= 8'b01000000;
mem[771] <= 8'b00100101;


// and $t0 $t0 $t2
mem[772] <= 8'b00001101;
mem[773] <= 8'b00001010;
mem[774] <= 8'b01000000;
mem[775] <= 8'b00010100;
//test 2
// addi $t0 $0 5
mem[808] <= 8'b00100100;
mem[809] <= 8'b00001000;
mem[810] <= 8'b00000000;
mem[811] <= 8'b00000101;

// add $t0 $t0 $s1
mem[812] <= 8'b00001101;
mem[813] <= 8'b00010011;
mem[814] <= 8'b01000000;
mem[815] <= 8'b00100000;

// addi $t0 $t0 7
mem[816] <= 8'b00100101;
mem[817] <= 8'b00001000;
mem[818] <= 8'b00000000;
mem[819] <= 8'b00000111;	

// lw $t0 0($0)
mem[900] <= 8'b01001000;
mem[901] <= 8'b00001000;
mem[902] <= 8'b00000000;
mem[903] <= 8'b00000000;
// addi $t0 $t0 7
mem[904] <= 8'b00100101;
mem[905] <= 8'b00001000;
mem[906] <= 8'b00000000;
mem[907] <= 8'b00000111;
// lw $t0 0($0)
mem[908] <= 8'b01001000;
mem[909] <= 8'b00001000;
mem[910] <= 8'b00000000;
mem[911] <= 8'b00000000;						
	end	 
   assign instruction = {mem[PC],mem[PC+1],mem[PC+2],mem[PC+3]}; 
endmodule