//declares a 32x32 register file.
module registerFile();
	
	// this module is not complete ... you should use these names to declare the register file unit 
	
	
reg [31:0] registers_i[31:0];
	
reg [31:0] registers_f[31:0];
	
endmodule