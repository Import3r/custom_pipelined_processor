module MA(op1,op2,op3,result,status);
input [7:0] op1,op2,op3;
output [7:0] result;
output reg [3:0] status;
wire [7:0] multiTemp;
wire [3:0] Stemp;
multi m1(op1,op2,multiTemp);
BAdder b1(multiTemp,op3,0,result,Stemp);
always@* begin
status[2] = Stemp[2];
end
endmodule
